// computer.v
module computer(clk, alu_result_out_bus);
  input clk;
  output [7:0] alu_result_out_bus;
  
  // cables relacionados al modulo de status
  wire [3:0] alu_flags_out_bus; // flags salientes de ALU
  wire [3:0] status_out_bus;    // flags salientes de Status
  
  // Recomiendo pasar todas estas señales para afuera para poder ser vistas en el waveform
  wire [7:0]    pc_out_bus;
  wire [7:0]    dm_out_bus;
  wire [14:0]   im_out_bus;
  
  wire [7:0]    regA_out_bus;
  wire [7:0]    regB_out_bus;
  wire [7:0]    muxA_out_bus;
  wire [7:0]    muxB_out_bus;
  wire [7:0]    mux_data_out_bus;
  
  // señales de control output-eadas por el control unit
  wire          L_PC_sig, D_W_sig, SD_sig; // load de PC, write enable a Data Memory, y selector de MUX data
  wire          LA_sig, LB_sig;            // loads de A y B 
  wire [1:0]    SB_sig, SA_sig;            // selectores de MUXs A y B
  wire [2:0]    S_alu_sig;                 // selector de la ALU

  // cables adicionales de numeros 0 y 1 para MUXs de A y B
  wire [7:0]    const0 = 8'b00000000;
  wire [7:0]    const1 = 8'b00000001;

  // slice de out bus de Instruction Memory para separar opcode y literal
  wire [6:0]    opcode = im_out_bus[14:8]; // 7 MSBs del instruction memory
  wire [7:0]    k8     = im_out_bus[7:0];  // literal; 8 LSBs del instruction memory


  /*======= CABLEADO DE MODULOS =======*/
  control_unit CU(
    .opcode(opcode),
    .flags_status(status_out_bus),
    .L_PC(L_PC_sig),
    .D_W(D_W_sig),
    .SD(SD_sig),
    .LA(LA_sig),
    .LB(LB_sig),
    .SA(SA_sig),
    .SB(SB_sig),
    .S_alu(S_alu_sig)
  );

  pc PC(
    .clk(clk),
    .pc(pc_out_bus)
  );

  instruction_memory IM(
    .address(pc_out_bus),
    .out(im_out_bus)
  );

  register regA(
    .clk(clk), 
    .data(alu_result_out_bus), 
    .load(LA_sig), 
    .out(regA_out_bus)
  );
  
  register regB(
    .clk(clk), 
    .data(alu_result_out_bus), 
    .load(LB_sig), 
    .out(regB_out_bus)
  );

  mux4 muxA(
    .e0(regA_out_bus), 
    .e1(regB_out_bus),
    .e2(const1),
    .e3(const0),
    .sel(SA_sig),
    .out(muxA_out_bus)
  );

  mux4 muxB(
    .e0(regB_out_bus), 
    .e1(dm_out_bus),
    .e2(k8),
    .e3(const0),
    .sel(SB_sig),
    .out(muxB_out_bus)
  );

  mux2 mux_data(
    .e0(k8),
    .e1(regB_out_bus),
    .s(SD_sig),
    .out(mux_data_out_bus)
  );

  data_memory DM(
    .clk(clk),
    .data_in(alu_result_out_bus),
    .address(mux_data_out_bus),
    .w(D_W_sig),
    .data_out(dm_out_bus)
  );

  alu ALU(
    .a(muxA_out_bus),
    .b(muxB_out_bus),
    .s(S_alu_sig),
    .result_out(alu_result_out_bus),
    .flags_out(alu_flags_out_bus)
  );

  status Status(
    .clk(clk),
    .flags_in(alu_flags_out_bus),
    .flags_out(status_out_bus)
  );

endmodule
